--Scrap File Data Path
